// megafunction wizard: %Pixel Buffer DMA Controller v13.0%
// GENERATION: XML
// DMA.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module DMA (
		input  wire        clk,                  //             clock_reset.clk
		input  wire        reset,                //       clock_reset_reset.reset
		input  wire        master_readdatavalid, // avalon_pixel_dma_master.readdatavalid
		input  wire        master_waitrequest,   //                        .waitrequest
		output wire [31:0] master_address,       //                        .address
		output wire        master_arbiterlock,   //                        .lock
		output wire        master_read,          //                        .read
		input  wire [31:0] master_readdata,      //                        .readdata
		input  wire [1:0]  slave_address,        //    avalon_control_slave.address
		input  wire [3:0]  slave_byteenable,     //                        .byteenable
		input  wire        slave_read,           //                        .read
		input  wire        slave_write,          //                        .write
		input  wire [31:0] slave_writedata,      //                        .writedata
		output wire [31:0] slave_readdata,       //                        .readdata
		input  wire        stream_ready,         //     avalon_pixel_source.ready
		output wire        stream_startofpacket, //                        .startofpacket
		output wire        stream_endofpacket,   //                        .endofpacket
		output wire        stream_valid,         //                        .valid
		output wire [29:0] stream_data           //                        .data
	);

	DMA_0002 dma_inst (
		.clk                  (clk),                  //             clock_reset.clk
		.reset                (reset),                //       clock_reset_reset.reset
		.master_readdatavalid (master_readdatavalid), // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (master_waitrequest),   //                        .waitrequest
		.master_address       (master_address),       //                        .address
		.master_arbiterlock   (master_arbiterlock),   //                        .lock
		.master_read          (master_read),          //                        .read
		.master_readdata      (master_readdata),      //                        .readdata
		.slave_address        (slave_address),        //    avalon_control_slave.address
		.slave_byteenable     (slave_byteenable),     //                        .byteenable
		.slave_read           (slave_read),           //                        .read
		.slave_write          (slave_write),          //                        .write
		.slave_writedata      (slave_writedata),      //                        .writedata
		.slave_readdata       (slave_readdata),       //                        .readdata
		.stream_ready         (stream_ready),         //     avalon_pixel_source.ready
		.stream_startofpacket (stream_startofpacket), //                        .startofpacket
		.stream_endofpacket   (stream_endofpacket),   //                        .endofpacket
		.stream_valid         (stream_valid),         //                        .valid
		.stream_data          (stream_data)           //                        .data
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2017 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_up_avalon_video_pixel_buffer_dma" version="13.0" >
// Retrieval info: 	<generic name="addr_mode" value="X-Y" />
// Retrieval info: 	<generic name="start_address" value="0" />
// Retrieval info: 	<generic name="back_start_address" value="0" />
// Retrieval info: 	<generic name="image_width" value="640" />
// Retrieval info: 	<generic name="image_height" value="480" />
// Retrieval info: 	<generic name="color_space" value="30-bit RGB" />
// Retrieval info: 	<generic name="AUTO_DEVICE_FAMILY" value="Cyclone IV E" />
// Retrieval info: 	<generic name="AUTO_CLOCK_RESET_CLOCK_RATE" value="-1" />
// Retrieval info: </instance>
// IPFS_FILES : DMA.vo
// RELATED_FILES: DMA.v, DMA_0002.v
